module sevenSegDigit (
input logic [3:0] digit,
output logic [6:0] displayBits
);


endmodule